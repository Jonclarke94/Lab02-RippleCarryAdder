//=========================================================================
// Name & Email must be EXACTLY as in Gradescope roster!
// Name: Jonathan Clarke
// Email: jclar084@ucr.edu
// 
// Assignment name: Lab02
// Lab section: 021
// TA: 
// 
// I hereby certify that I have not received assistance on this assignment,
// or used code, from ANY outside source other than the instruction team
// (apart from what was provided in the starter file).
//
//=========================================================================

`timescale 1ns / 1ps

//  Constant definitions 

module ripple_carry_adder # ( parameter NUMBITS = 16 ) (
    input  wire[NUMBITS-1:0] A, 
    input  wire[NUMBITS-1:0] B, 
    input wire carryin, 
    output reg [NUMBITS-1:0] result,  
    output reg carryout); 

    // ------------------------------
    // Insert your solution below
    // ------------------------------ 
     reg carry;

    always @* begin
        carry = carryin;
        result = 0;
        for (int i=0; i<NUMBITS; i=i+1) begin
            result[i] = A[i] ^ B[i] ^ carry;
            carry = (A[i] & B[i]) | (carry & (A[i] ^ B[i]));
        end
        carryout = carry;
    end

endmodule
